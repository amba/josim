
* DC_SFQ converter
* NEW RSFQ CIRCUITS S.V. Polonsky et al.
* See Fig 3a

.subckt DC_SFQ 10
.param tstep=100p

.param idc_in=500u
IDC    0          1          pwl(0    0  tstep  idc_in 2*tstep idc_in 3*tstep 0 4*tstep 0 5*tstep idc_in 6*tstep idc_in 7*tstep 0 8*tstep 0 9*tstep idc_in 10*tstep idc_in 11*tstep 0 12*tstep 0 13*tstep idc_in 14*tstep idc_in 15*tstep 0 16*tstep 0)
IBIAS1   0         5          pwl(0 0 5p 400u)
IBIAS2   0         8          pwl(0 0 5p 380u)
B1      3         4           jjmod
B2      2         4           jjmod
B3      4         0           jjmod
B4      6         0           jjmod
B5      7         0           jjmod
B6      9         0           jjmod
L1      1         3           1.4p
L2      1         2           1.3p
L3      2         0           2.5p
L4      4         5           0.4p
L5      5         6           1.2p
L6      6         7           2.4p
L7      7         8           2p
L8      8         9           2p
L9      9         10          4p
.model jjmod jj(rtype=1, vg=2mV, cap=1fF, r0=10, rN=10, icrit=250uA)
.ends

.subckt SPLITTER 1 7 10
L2 5 7      1p
L3 5 10      1p
L4 1 2      1p
L5 2 3      1p
L6 3 4      1p
L7 4 5      1p
B1 7 0          jjmod    area=2.5
B2 10 0		jjmod    area=2.5
B5 2 0		jjmod    area=2.5
B6 4 0		jjmod    area=2.5
I1   0         3          pwl(0 0 1p 450u)
.model jjmod jj(rtype=1, vg=2mV, cap=1fF, r0=10, rN=10, icrit=100uA)
.ends


.subckt TFLIPFLOP 1 8 11
L1 7 10     8p
L2 5 6      0.14p
L3 5 9      1.87p
L4 1 2      2.67p
L5 2 3      1.33p
L6 3 4      0.8p
L7 4 5      0.27p
L8 7 8      8p
L12 10 11   5.33p
B1 7 0          jjmod    area=1.25
B2 10 0		jjmod    area=1.92
B3 6 7		jjmod    area=3
B4 9 10		jjmod    area=1.25
B5 2 0		jjmod    area=2.5
B6 4 0		jjmod    area=2.5
B7 8 0		jjmod    area=1.25
B9 11 0         jjmod    area=1.92
I1   0         3          pwl(0 0 1p 450u)
.model jjmod jj(rtype=1, vg=2mV, cap=1fF, r0=10, rN=10, icrit=100uA)
.ends


XIN DC_SFQ 1
XS SPLITTER 1 2 3
* XT TFLIPFLOP 1 2 3
ROUT1 2 0 100
ROUT2 3 0 100
.tran 0.1p 2000p 0 0.1p
.print DEVI IDC.XIN
.print PHASE B6.XS
.print PHASE B1.XS
.print PHASE 1
.print DEVI ROUT1
.print DEVI ROUT2
