.param vdc_in=0.1
.param tstep=10000p
.param deltat=0.01p

VDC    0          1          pwl(0    0  tstep  vdc_in)
R1     1          2          300
R2     3          2          300
VAC    0          3          sin(0    vdc_in*1 200e9)
B1      2         0           jjmod

.model jjmod jj(rtype=1, vg=2.8e-3, cap=10fF, r0=100, rN=25, icrit=0.2e-3)

.tran deltat tstep
.print DEVI B1
.print DEVV B1
# .print PHASE B1
